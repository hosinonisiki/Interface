LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.Numeric_std.ALL;

ENTITY WaveGen IS
    PORT(
        
    );
END WaveGen;