LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.Numeric_std.ALL;

ENTITY FIR_10M IS
    PORT(
        SIGNAL input : IN signed(15 DOWNTO 0);
        SIGNAL output : OUT signed(15 DOWNTO 0);
        SIGNAL Reset : IN std_logic;
        SIGNAL Clk : IN std_logic
    );
END FIR_10M;

ARCHITECTURE bhvr OF FIR_10M IS
    CONSTANT tap : INTEGER := 256;
    TYPE envelope_array IS ARRAY(0 TO 255) OF signed(11 DOWNTO 0);
    CONSTANT LUT_envelope : envelope_array := (
        "000000000000",
        "111111110000",
        "111111100001",
        "111111010010",
        "111111000101",
        "111110111010",
        "111110110010",
        "111110101100",
        "111110101010",
        "111110101011",
        "111110101111",
        "111110110110",
        "111111000001",
        "111111001110",
        "111111011110",
        "111111101111",
        "000000000000",
        "000000010010",
        "000000100100",
        "000000110101",
        "000001000100",
        "000001010001",
        "000001011010",
        "000001100001",
        "000001100100",
        "000001100011",
        "000001011110",
        "000001010101",
        "000001001001",
        "000000111010",
        "000000101000",
        "000000010100",
        "000000000000",
        "111111101011",
        "111111010110",
        "111111000010",
        "111110110000",
        "111110100001",
        "111110010101",
        "111110001110",
        "111110001010",
        "111110001011",
        "111110010001",
        "111110011011",
        "111110101001",
        "111110111011",
        "111111010000",
        "111111100111",
        "000000000000",
        "000000011001",
        "000000110011",
        "000001001011",
        "000001100000",
        "000001110011",
        "000010000010",
        "000010001100",
        "000010010000",
        "000010010000",
        "000010001001",
        "000001111101",
        "000001101100",
        "000001010110",
        "000000111100",
        "000000011111",
        "000000000000",
        "111111100000",
        "111111000000",
        "111110100010",
        "111110000110",
        "111101101110",
        "111101011010",
        "111101001101",
        "111101000110",
        "111101000111",
        "111101001110",
        "111101011101",
        "111101110011",
        "111110001111",
        "111110110001",
        "111111010111",
        "000000000000",
        "000000101011",
        "000001010110",
        "000010000000",
        "000010100111",
        "000011001001",
        "000011100101",
        "000011111001",
        "000100000100",
        "000100000110",
        "000011111101",
        "000011101010",
        "000011001100",
        "000010100101",
        "000001110101",
        "000000111101",
        "000000000000",
        "111110111111",
        "111101111100",
        "111100111001",
        "111011111001",
        "111010111111",
        "111010001110",
        "111001101000",
        "111001001110",
        "111001000100",
        "111001001011",
        "111001100100",
        "111010010000",
        "111011010000",
        "111100100011",
        "111110001001",
        "000000000000",
        "000010000111",
        "000100011100",
        "000110111101",
        "001001100110",
        "001100010100",
        "001111000011",
        "010001110000",
        "010100010111",
        "010110110100",
        "011001000101",
        "011011000101",
        "011100110010",
        "011110001010",
        "011111001010",
        "011111110001",
        "011111111111",
        "011111110001",
        "011111001010",
        "011110001010",
        "011100110010",
        "011011000101",
        "011001000101",
        "010110110100",
        "010100010111",
        "010001110000",
        "001111000011",
        "001100010100",
        "001001100110",
        "000110111101",
        "000100011100",
        "000010000111",
        "000000000000",
        "111110001001",
        "111100100011",
        "111011010000",
        "111010010000",
        "111001100100",
        "111001001011",
        "111001000100",
        "111001001110",
        "111001101000",
        "111010001110",
        "111010111111",
        "111011111001",
        "111100111001",
        "111101111100",
        "111110111111",
        "000000000000",
        "000000111101",
        "000001110101",
        "000010100101",
        "000011001100",
        "000011101010",
        "000011111101",
        "000100000110",
        "000100000100",
        "000011111001",
        "000011100101",
        "000011001001",
        "000010100111",
        "000010000000",
        "000001010110",
        "000000101011",
        "000000000000",
        "111111010111",
        "111110110001",
        "111110001111",
        "111101110011",
        "111101011101",
        "111101001110",
        "111101000111",
        "111101000110",
        "111101001101",
        "111101011010",
        "111101101110",
        "111110000110",
        "111110100010",
        "111111000000",
        "111111100000",
        "000000000000",
        "000000011111",
        "000000111100",
        "000001010110",
        "000001101100",
        "000001111101",
        "000010001001",
        "000010010000",
        "000010010000",
        "000010001100",
        "000010000010",
        "000001110011",
        "000001100000",
        "000001001011",
        "000000110011",
        "000000011001",
        "000000000000",
        "111111100111",
        "111111010000",
        "111110111011",
        "111110101001",
        "111110011011",
        "111110010001",
        "111110001011",
        "111110001010",
        "111110001110",
        "111110010101",
        "111110100001",
        "111110110000",
        "111111000010",
        "111111010110",
        "111111101011",
        "000000000000",
        "000000010100",
        "000000101000",
        "000000111010",
        "000001001001",
        "000001010101",
        "000001011110",
        "000001100011",
        "000001100100",
        "000001100001",
        "000001011010",
        "000001010001",
        "000001000100",
        "000000110101",
        "000000100100",
        "000000010010",
        "000000000000",
        "111111101111",
        "111111011110",
        "111111001110",
        "111111000001",
        "111110110110",
        "111110101111",
        "111110101011",
        "111110101010",
        "111110101100",
        "111110110010",
        "111110111010",
        "111111000101",
        "111111010010",
        "111111100001",
        "111111110000"     
    );
    TYPE source_array IS ARRAY(0 TO 255) OF signed(15 DOWNTO 0);
    SIGNAL source : source_array;
    TYPE image_array IS ARRAY(0 TO 255) OF signed(27 DOWNTO 0);
    SIGNAL image : image_array;
    TYPE sum_array IS ARRAY(0 TO 254) OF signed(19 DOWNTO 0);
    SIGNAL sum : sum_array;
    TYPE constant_array IS ARRAY(0 TO 7) OF INTEGER;
    CONSTANT adders_per_row : constant_array := (
        128, 64, 32, 16, 8, 4, 2, 1
    );
    CONSTANT adders_starting_number : constant_array := (
        0, 128, 192, 224, 240, 248, 252, 254
    );
BEGIN
    PROCESS(Clk)
    BEGIN
        IF rising_edge(Clk) THEN
            source(0) <= input;
            output <= sum(254)(19 DOWNTO 4);
        END IF;
    END PROCESS;
    image(0) <= source(0) * LUT_envelope(0);
    gen_multiplication : FOR i IN 0 TO 254 GENERATE
        PROCESS(Clk)
        BEGIN
            IF rising_edge(Clk) THEN
                source(i + 1) <= source(i);
            END IF;
        END PROCESS;
        image(i + 1) <= source(i + 1) * LUT_envelope(i + 1);
        gen_sum_first_row : IF (i MOD 2 = 0) GENERATE
            PROCESS(Clk)
            BEGIN
                IF rising_edge(Clk) THEN
                    sum(i / 2) <= ((7 DOWNTO 0 => image(i)(27)) & image(i)(27 DOWNTO 16)) + ((7 DOWNTO 0 => image(i + 1)(27)) & image(i + 1)(27 DOWNTO 16));
                END IF;
            END PROCESS;
        END GENERATE gen_sum_first_row; 
    END GENERATE gen_multiplication;
-- 0 1 2 3 4 5 6 7
--  8   9  10  11
--    12    13
--       14
    gen_sum_row : FOR i IN 0 TO 6 GENERATE
        gen_sum : FOR j IN 0 TO adders_per_row(i + 1) - 1 GENERATE
            PROCESS(Clk)
            BEGIN
                IF rising_edge(Clk) THEN
                    sum(j + adders_starting_number(i + 1)) <= sum(j * 2 + adders_starting_number(i)) + sum(j * 2 + adders_starting_number(i) + 1);
                END IF;
            END PROCESS;
        END GENERATE gen_sum;
    END GENERATE gen_sum_row;
END bhvr;